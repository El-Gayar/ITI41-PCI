`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:20:59 02/16/2021 
// Design Name: 
// Module Name:    add_data 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module add_data(
    input clk,
    input rst,
    inout [31:0] ad,
	 inout [3:0]  c_be,
	 inout par,
    );


endmodule
